module counterDebouncer #(parameter C_MAX = 500000)(
	input clk, rst_a,
	output reg flag_check
);

reg[18:0] counter_reg_aux;

always @(posedge clk or negedge rst_a)
begin
	if(!rst_a) //if(rst_a == 0) si el reset es igual a 0
	begin
		counter_reg_aux <= 0;
		flag_check  <= 0;
	end
	else
	begin
		if(counter_reg_aux >= C_MAX)
		begin
			counter_reg_aux <= 0;
			flag_check <= 1;
		end
		else
		begin
			counter_reg_aux <= counter_reg_aux + 1;
			flag_check <= 0;
		end
	end

end
endmodule